library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
entity Comparator_2_Digit_TB is

end Comparator_2_Digit_TB;

architecture Behavioral of Comparator_2_Digit_TB is
component Comparator_2_Digit
begin


end Behavioral;
