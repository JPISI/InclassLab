library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity Full_adder_structural_TB is
end Full_adder_structural_TB;

architecture Behavioral of Full_adder_structural_TB is
  signal A, B, Cin, S, Cout : std_logic;
  
  uut: entity Full_adder_structural
  port map
begin


end Behavioral;
